`timescale 1 ns/100 ps
// Version: PolarFire v2.2 12.200.30.10


module Init_Monitor_Init_Monitor_0_PF_INIT_MONITOR(
       FABRIC_POR_N,
       PCIE_INIT_DONE,
       SRAM_INIT_DONE,
       DEVICE_INIT_DONE,
       USRAM_INIT_DONE,
       XCVR_INIT_DONE,
       USRAM_INIT_FROM_SNVM_DONE,
       USRAM_INIT_FROM_UPROM_DONE,
       USRAM_INIT_FROM_SPI_DONE,
       SRAM_INIT_FROM_SNVM_DONE,
       SRAM_INIT_FROM_UPROM_DONE,
       SRAM_INIT_FROM_SPI_DONE,
       AUTOCALIB_DONE
    );
output FABRIC_POR_N;
output PCIE_INIT_DONE;
output SRAM_INIT_DONE;
output DEVICE_INIT_DONE;
output USRAM_INIT_DONE;
output XCVR_INIT_DONE;
output USRAM_INIT_FROM_SNVM_DONE;
output USRAM_INIT_FROM_UPROM_DONE;
output USRAM_INIT_FROM_SPI_DONE;
output SRAM_INIT_FROM_SNVM_DONE;
output SRAM_INIT_FROM_UPROM_DONE;
output SRAM_INIT_FROM_SPI_DONE;
output AUTOCALIB_DONE;

    wire GND_net, VCC_net;
    
    INIT #( .FABRIC_POR_N_SIMULATION_DELAY(1000), .PCIE_INIT_DONE_SIMULATION_DELAY(4000)
        , .SRAM_INIT_DONE_SIMULATION_DELAY(6000), .UIC_INIT_DONE_SIMULATION_DELAY(7000)
        , .USRAM_INIT_DONE_SIMULATION_DELAY(5000) )  I_INIT (
        .FABRIC_POR_N(FABRIC_POR_N), .GPIO_ACTIVE(), .HSIO_ACTIVE(), 
        .PCIE_INIT_DONE(PCIE_INIT_DONE), .RFU({AUTOCALIB_DONE, nc0, 
        nc1, nc2, nc3, SRAM_INIT_FROM_SPI_DONE, 
        SRAM_INIT_FROM_UPROM_DONE, SRAM_INIT_FROM_SNVM_DONE, 
        USRAM_INIT_FROM_SPI_DONE, USRAM_INIT_FROM_UPROM_DONE, 
        USRAM_INIT_FROM_SNVM_DONE, XCVR_INIT_DONE}), .SRAM_INIT_DONE(
        SRAM_INIT_DONE), .UIC_INIT_DONE(DEVICE_INIT_DONE), 
        .USRAM_INIT_DONE(USRAM_INIT_DONE));
    VCC vcc_inst (.Y(VCC_net));
    GND gnd_inst (.Y(GND_net));
    
endmodule
