`timescale 1 ns/100 ps
// Version: PolarFire v2.2 12.200.30.10


module LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM(
       W_DATA,
       R_DATA,
       W_ADDR,
       R_ADDR,
       W_EN,
       R_EN,
       CLK,
       WBYTE_EN
    );
input  [39:0] W_DATA;
output [39:0] R_DATA;
input  [13:0] W_ADDR;
input  [13:0] R_ADDR;
input  W_EN;
input  R_EN;
input  CLK;
input  [39:0] WBYTE_EN;

    wire \ACCESS_BUSY[0][0] , \SB_CORRECT[0][0] , \DB_DETECT[0][0] , 
        \ACCESS_BUSY[0][1] , \SB_CORRECT[0][1] , \DB_DETECT[0][1] , 
        \ACCESS_BUSY[0][2] , \SB_CORRECT[0][2] , \DB_DETECT[0][2] , 
        \ACCESS_BUSY[0][3] , \SB_CORRECT[0][3] , \DB_DETECT[0][3] , 
        \ACCESS_BUSY[0][4] , \SB_CORRECT[0][4] , \DB_DETECT[0][4] , 
        \ACCESS_BUSY[0][5] , \SB_CORRECT[0][5] , \DB_DETECT[0][5] , 
        \ACCESS_BUSY[0][6] , \SB_CORRECT[0][6] , \DB_DETECT[0][6] , 
        \ACCESS_BUSY[0][7] , \SB_CORRECT[0][7] , \DB_DETECT[0][7] , 
        \ACCESS_BUSY[0][8] , \SB_CORRECT[0][8] , \DB_DETECT[0][8] , 
        \ACCESS_BUSY[0][9] , \SB_CORRECT[0][9] , \DB_DETECT[0][9] , 
        \ACCESS_BUSY[0][10] , \SB_CORRECT[0][10] , \DB_DETECT[0][10] , 
        \ACCESS_BUSY[0][11] , \SB_CORRECT[0][11] , \DB_DETECT[0][11] , 
        \ACCESS_BUSY[0][12] , \SB_CORRECT[0][12] , \DB_DETECT[0][12] , 
        \ACCESS_BUSY[0][13] , \SB_CORRECT[0][13] , \DB_DETECT[0][13] , 
        \ACCESS_BUSY[0][14] , \SB_CORRECT[0][14] , \DB_DETECT[0][14] , 
        \ACCESS_BUSY[0][15] , \SB_CORRECT[0][15] , \DB_DETECT[0][15] , 
        \ACCESS_BUSY[0][16] , \SB_CORRECT[0][16] , \DB_DETECT[0][16] , 
        \ACCESS_BUSY[0][17] , \SB_CORRECT[0][17] , \DB_DETECT[0][17] , 
        \ACCESS_BUSY[0][18] , \SB_CORRECT[0][18] , \DB_DETECT[0][18] , 
        \ACCESS_BUSY[0][19] , \SB_CORRECT[0][19] , \DB_DETECT[0][19] , 
        \ACCESS_BUSY[0][20] , \SB_CORRECT[0][20] , \DB_DETECT[0][20] , 
        \ACCESS_BUSY[0][21] , \SB_CORRECT[0][21] , \DB_DETECT[0][21] , 
        \ACCESS_BUSY[0][22] , \SB_CORRECT[0][22] , \DB_DETECT[0][22] , 
        \ACCESS_BUSY[0][23] , \SB_CORRECT[0][23] , \DB_DETECT[0][23] , 
        \ACCESS_BUSY[0][24] , \SB_CORRECT[0][24] , \DB_DETECT[0][24] , 
        \ACCESS_BUSY[0][25] , \SB_CORRECT[0][25] , \DB_DETECT[0][25] , 
        \ACCESS_BUSY[0][26] , \SB_CORRECT[0][26] , \DB_DETECT[0][26] , 
        \ACCESS_BUSY[0][27] , \SB_CORRECT[0][27] , \DB_DETECT[0][27] , 
        \ACCESS_BUSY[0][28] , \SB_CORRECT[0][28] , \DB_DETECT[0][28] , 
        \ACCESS_BUSY[0][29] , \SB_CORRECT[0][29] , \DB_DETECT[0][29] , 
        \ACCESS_BUSY[0][30] , \SB_CORRECT[0][30] , \DB_DETECT[0][30] , 
        \ACCESS_BUSY[0][31] , \SB_CORRECT[0][31] , \DB_DETECT[0][31] , 
        \ACCESS_BUSY[0][32] , \SB_CORRECT[0][32] , \DB_DETECT[0][32] , 
        \ACCESS_BUSY[0][33] , \SB_CORRECT[0][33] , \DB_DETECT[0][33] , 
        \ACCESS_BUSY[0][34] , \SB_CORRECT[0][34] , \DB_DETECT[0][34] , 
        \ACCESS_BUSY[0][35] , \SB_CORRECT[0][35] , \DB_DETECT[0][35] , 
        \ACCESS_BUSY[0][36] , \SB_CORRECT[0][36] , \DB_DETECT[0][36] , 
        \ACCESS_BUSY[0][37] , \SB_CORRECT[0][37] , \DB_DETECT[0][37] , 
        \ACCESS_BUSY[0][38] , \SB_CORRECT[0][38] , \DB_DETECT[0][38] , 
        \ACCESS_BUSY[0][39] , \SB_CORRECT[0][39] , \DB_DETECT[0][39] , 
        VCC, GND, ADLIB_VCC;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign ADLIB_VCC = VCC_power_net1;
    
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%34%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C34 (.A_DOUT({
        nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7, nc8, nc9, nc10, nc11, 
        nc12, nc13, nc14, nc15, nc16, nc17, nc18, R_DATA[34]}), 
        .B_DOUT({nc19, nc20, nc21, nc22, nc23, nc24, nc25, nc26, nc27, 
        nc28, nc29, nc30, nc31, nc32, nc33, nc34, nc35, nc36, nc37, 
        nc38}), .DB_DETECT(\DB_DETECT[0][34] ), .SB_CORRECT(
        \SB_CORRECT[0][34] ), .ACCESS_BUSY(\ACCESS_BUSY[0][34] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[34]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[34]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%24%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C24 (.A_DOUT({
        nc39, nc40, nc41, nc42, nc43, nc44, nc45, nc46, nc47, nc48, 
        nc49, nc50, nc51, nc52, nc53, nc54, nc55, nc56, nc57, 
        R_DATA[24]}), .B_DOUT({nc58, nc59, nc60, nc61, nc62, nc63, 
        nc64, nc65, nc66, nc67, nc68, nc69, nc70, nc71, nc72, nc73, 
        nc74, nc75, nc76, nc77}), .DB_DETECT(\DB_DETECT[0][24] ), 
        .SB_CORRECT(\SB_CORRECT[0][24] ), .ACCESS_BUSY(
        \ACCESS_BUSY[0][24] ), .A_ADDR({R_ADDR[13], R_ADDR[12], 
        R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK)
        , .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), .A_REN(
        R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC)
        , .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], W_ADDR[12], 
        W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], W_ADDR[7], 
        W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], W_ADDR[2], 
        W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, W_DATA[24]}), 
        .B_REN(VCC), .B_WEN({GND, WBYTE_EN[24]}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), 
        .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%31%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C31 (.A_DOUT({
        nc78, nc79, nc80, nc81, nc82, nc83, nc84, nc85, nc86, nc87, 
        nc88, nc89, nc90, nc91, nc92, nc93, nc94, nc95, nc96, 
        R_DATA[31]}), .B_DOUT({nc97, nc98, nc99, nc100, nc101, nc102, 
        nc103, nc104, nc105, nc106, nc107, nc108, nc109, nc110, nc111, 
        nc112, nc113, nc114, nc115, nc116}), .DB_DETECT(
        \DB_DETECT[0][31] ), .SB_CORRECT(\SB_CORRECT[0][31] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][31] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[31]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[31]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%32%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C32 (.A_DOUT({
        nc117, nc118, nc119, nc120, nc121, nc122, nc123, nc124, nc125, 
        nc126, nc127, nc128, nc129, nc130, nc131, nc132, nc133, nc134, 
        nc135, R_DATA[32]}), .B_DOUT({nc136, nc137, nc138, nc139, 
        nc140, nc141, nc142, nc143, nc144, nc145, nc146, nc147, nc148, 
        nc149, nc150, nc151, nc152, nc153, nc154, nc155}), .DB_DETECT(
        \DB_DETECT[0][32] ), .SB_CORRECT(\SB_CORRECT[0][32] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][32] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[32]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[32]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%33%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C33 (.A_DOUT({
        nc156, nc157, nc158, nc159, nc160, nc161, nc162, nc163, nc164, 
        nc165, nc166, nc167, nc168, nc169, nc170, nc171, nc172, nc173, 
        nc174, R_DATA[33]}), .B_DOUT({nc175, nc176, nc177, nc178, 
        nc179, nc180, nc181, nc182, nc183, nc184, nc185, nc186, nc187, 
        nc188, nc189, nc190, nc191, nc192, nc193, nc194}), .DB_DETECT(
        \DB_DETECT[0][33] ), .SB_CORRECT(\SB_CORRECT[0][33] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][33] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[33]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[33]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%22%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C22 (.A_DOUT({
        nc195, nc196, nc197, nc198, nc199, nc200, nc201, nc202, nc203, 
        nc204, nc205, nc206, nc207, nc208, nc209, nc210, nc211, nc212, 
        nc213, R_DATA[22]}), .B_DOUT({nc214, nc215, nc216, nc217, 
        nc218, nc219, nc220, nc221, nc222, nc223, nc224, nc225, nc226, 
        nc227, nc228, nc229, nc230, nc231, nc232, nc233}), .DB_DETECT(
        \DB_DETECT[0][22] ), .SB_CORRECT(\SB_CORRECT[0][22] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][22] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[22]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[22]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%23%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C23 (.A_DOUT({
        nc234, nc235, nc236, nc237, nc238, nc239, nc240, nc241, nc242, 
        nc243, nc244, nc245, nc246, nc247, nc248, nc249, nc250, nc251, 
        nc252, R_DATA[23]}), .B_DOUT({nc253, nc254, nc255, nc256, 
        nc257, nc258, nc259, nc260, nc261, nc262, nc263, nc264, nc265, 
        nc266, nc267, nc268, nc269, nc270, nc271, nc272}), .DB_DETECT(
        \DB_DETECT[0][23] ), .SB_CORRECT(\SB_CORRECT[0][23] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][23] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[23]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[23]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%21%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C21 (.A_DOUT({
        nc273, nc274, nc275, nc276, nc277, nc278, nc279, nc280, nc281, 
        nc282, nc283, nc284, nc285, nc286, nc287, nc288, nc289, nc290, 
        nc291, R_DATA[21]}), .B_DOUT({nc292, nc293, nc294, nc295, 
        nc296, nc297, nc298, nc299, nc300, nc301, nc302, nc303, nc304, 
        nc305, nc306, nc307, nc308, nc309, nc310, nc311}), .DB_DETECT(
        \DB_DETECT[0][21] ), .SB_CORRECT(\SB_CORRECT[0][21] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][21] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[21]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[21]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%9%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C9 (.A_DOUT({
        nc312, nc313, nc314, nc315, nc316, nc317, nc318, nc319, nc320, 
        nc321, nc322, nc323, nc324, nc325, nc326, nc327, nc328, nc329, 
        nc330, R_DATA[9]}), .B_DOUT({nc331, nc332, nc333, nc334, nc335, 
        nc336, nc337, nc338, nc339, nc340, nc341, nc342, nc343, nc344, 
        nc345, nc346, nc347, nc348, nc349, nc350}), .DB_DETECT(
        \DB_DETECT[0][9] ), .SB_CORRECT(\SB_CORRECT[0][9] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][9] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[9]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[9]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%19%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C19 (.A_DOUT({
        nc351, nc352, nc353, nc354, nc355, nc356, nc357, nc358, nc359, 
        nc360, nc361, nc362, nc363, nc364, nc365, nc366, nc367, nc368, 
        nc369, R_DATA[19]}), .B_DOUT({nc370, nc371, nc372, nc373, 
        nc374, nc375, nc376, nc377, nc378, nc379, nc380, nc381, nc382, 
        nc383, nc384, nc385, nc386, nc387, nc388, nc389}), .DB_DETECT(
        \DB_DETECT[0][19] ), .SB_CORRECT(\SB_CORRECT[0][19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][19] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[19]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[19]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%8%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C8 (.A_DOUT({
        nc390, nc391, nc392, nc393, nc394, nc395, nc396, nc397, nc398, 
        nc399, nc400, nc401, nc402, nc403, nc404, nc405, nc406, nc407, 
        nc408, R_DATA[8]}), .B_DOUT({nc409, nc410, nc411, nc412, nc413, 
        nc414, nc415, nc416, nc417, nc418, nc419, nc420, nc421, nc422, 
        nc423, nc424, nc425, nc426, nc427, nc428}), .DB_DETECT(
        \DB_DETECT[0][8] ), .SB_CORRECT(\SB_CORRECT[0][8] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][8] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[8]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[8]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%37%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C37 (.A_DOUT({
        nc429, nc430, nc431, nc432, nc433, nc434, nc435, nc436, nc437, 
        nc438, nc439, nc440, nc441, nc442, nc443, nc444, nc445, nc446, 
        nc447, R_DATA[37]}), .B_DOUT({nc448, nc449, nc450, nc451, 
        nc452, nc453, nc454, nc455, nc456, nc457, nc458, nc459, nc460, 
        nc461, nc462, nc463, nc464, nc465, nc466, nc467}), .DB_DETECT(
        \DB_DETECT[0][37] ), .SB_CORRECT(\SB_CORRECT[0][37] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][37] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[37]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[37]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%1%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C1 (.A_DOUT({
        nc468, nc469, nc470, nc471, nc472, nc473, nc474, nc475, nc476, 
        nc477, nc478, nc479, nc480, nc481, nc482, nc483, nc484, nc485, 
        nc486, R_DATA[1]}), .B_DOUT({nc487, nc488, nc489, nc490, nc491, 
        nc492, nc493, nc494, nc495, nc496, nc497, nc498, nc499, nc500, 
        nc501, nc502, nc503, nc504, nc505, nc506}), .DB_DETECT(
        \DB_DETECT[0][1] ), .SB_CORRECT(\SB_CORRECT[0][1] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][1] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[1]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[1]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%27%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C27 (.A_DOUT({
        nc507, nc508, nc509, nc510, nc511, nc512, nc513, nc514, nc515, 
        nc516, nc517, nc518, nc519, nc520, nc521, nc522, nc523, nc524, 
        nc525, R_DATA[27]}), .B_DOUT({nc526, nc527, nc528, nc529, 
        nc530, nc531, nc532, nc533, nc534, nc535, nc536, nc537, nc538, 
        nc539, nc540, nc541, nc542, nc543, nc544, nc545}), .DB_DETECT(
        \DB_DETECT[0][27] ), .SB_CORRECT(\SB_CORRECT[0][27] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][27] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[27]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[27]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%10%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C10 (.A_DOUT({
        nc546, nc547, nc548, nc549, nc550, nc551, nc552, nc553, nc554, 
        nc555, nc556, nc557, nc558, nc559, nc560, nc561, nc562, nc563, 
        nc564, R_DATA[10]}), .B_DOUT({nc565, nc566, nc567, nc568, 
        nc569, nc570, nc571, nc572, nc573, nc574, nc575, nc576, nc577, 
        nc578, nc579, nc580, nc581, nc582, nc583, nc584}), .DB_DETECT(
        \DB_DETECT[0][10] ), .SB_CORRECT(\SB_CORRECT[0][10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][10] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[10]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[10]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%4%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C4 (.A_DOUT({
        nc585, nc586, nc587, nc588, nc589, nc590, nc591, nc592, nc593, 
        nc594, nc595, nc596, nc597, nc598, nc599, nc600, nc601, nc602, 
        nc603, R_DATA[4]}), .B_DOUT({nc604, nc605, nc606, nc607, nc608, 
        nc609, nc610, nc611, nc612, nc613, nc614, nc615, nc616, nc617, 
        nc618, nc619, nc620, nc621, nc622, nc623}), .DB_DETECT(
        \DB_DETECT[0][4] ), .SB_CORRECT(\SB_CORRECT[0][4] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][4] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[4]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[4]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%16%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C16 (.A_DOUT({
        nc624, nc625, nc626, nc627, nc628, nc629, nc630, nc631, nc632, 
        nc633, nc634, nc635, nc636, nc637, nc638, nc639, nc640, nc641, 
        nc642, R_DATA[16]}), .B_DOUT({nc643, nc644, nc645, nc646, 
        nc647, nc648, nc649, nc650, nc651, nc652, nc653, nc654, nc655, 
        nc656, nc657, nc658, nc659, nc660, nc661, nc662}), .DB_DETECT(
        \DB_DETECT[0][16] ), .SB_CORRECT(\SB_CORRECT[0][16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][16] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[16]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[16]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%18%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C18 (.A_DOUT({
        nc663, nc664, nc665, nc666, nc667, nc668, nc669, nc670, nc671, 
        nc672, nc673, nc674, nc675, nc676, nc677, nc678, nc679, nc680, 
        nc681, R_DATA[18]}), .B_DOUT({nc682, nc683, nc684, nc685, 
        nc686, nc687, nc688, nc689, nc690, nc691, nc692, nc693, nc694, 
        nc695, nc696, nc697, nc698, nc699, nc700, nc701}), .DB_DETECT(
        \DB_DETECT[0][18] ), .SB_CORRECT(\SB_CORRECT[0][18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][18] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[18]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[18]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%0%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0 (.A_DOUT({
        nc702, nc703, nc704, nc705, nc706, nc707, nc708, nc709, nc710, 
        nc711, nc712, nc713, nc714, nc715, nc716, nc717, nc718, nc719, 
        nc720, R_DATA[0]}), .B_DOUT({nc721, nc722, nc723, nc724, nc725, 
        nc726, nc727, nc728, nc729, nc730, nc731, nc732, nc733, nc734, 
        nc735, nc736, nc737, nc738, nc739, nc740}), .DB_DETECT(
        \DB_DETECT[0][0] ), .SB_CORRECT(\SB_CORRECT[0][0] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][0] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%15%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C15 (.A_DOUT({
        nc741, nc742, nc743, nc744, nc745, nc746, nc747, nc748, nc749, 
        nc750, nc751, nc752, nc753, nc754, nc755, nc756, nc757, nc758, 
        nc759, R_DATA[15]}), .B_DOUT({nc760, nc761, nc762, nc763, 
        nc764, nc765, nc766, nc767, nc768, nc769, nc770, nc771, nc772, 
        nc773, nc774, nc775, nc776, nc777, nc778, nc779}), .DB_DETECT(
        \DB_DETECT[0][15] ), .SB_CORRECT(\SB_CORRECT[0][15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][15] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[15]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[15]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%5%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C5 (.A_DOUT({
        nc780, nc781, nc782, nc783, nc784, nc785, nc786, nc787, nc788, 
        nc789, nc790, nc791, nc792, nc793, nc794, nc795, nc796, nc797, 
        nc798, R_DATA[5]}), .B_DOUT({nc799, nc800, nc801, nc802, nc803, 
        nc804, nc805, nc806, nc807, nc808, nc809, nc810, nc811, nc812, 
        nc813, nc814, nc815, nc816, nc817, nc818}), .DB_DETECT(
        \DB_DETECT[0][5] ), .SB_CORRECT(\SB_CORRECT[0][5] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][5] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[5]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[5]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%39%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C39 (.A_DOUT({
        nc819, nc820, nc821, nc822, nc823, nc824, nc825, nc826, nc827, 
        nc828, nc829, nc830, nc831, nc832, nc833, nc834, nc835, nc836, 
        nc837, R_DATA[39]}), .B_DOUT({nc838, nc839, nc840, nc841, 
        nc842, nc843, nc844, nc845, nc846, nc847, nc848, nc849, nc850, 
        nc851, nc852, nc853, nc854, nc855, nc856, nc857}), .DB_DETECT(
        \DB_DETECT[0][39] ), .SB_CORRECT(\SB_CORRECT[0][39] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][39] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[39]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[39]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%29%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C29 (.A_DOUT({
        nc858, nc859, nc860, nc861, nc862, nc863, nc864, nc865, nc866, 
        nc867, nc868, nc869, nc870, nc871, nc872, nc873, nc874, nc875, 
        nc876, R_DATA[29]}), .B_DOUT({nc877, nc878, nc879, nc880, 
        nc881, nc882, nc883, nc884, nc885, nc886, nc887, nc888, nc889, 
        nc890, nc891, nc892, nc893, nc894, nc895, nc896}), .DB_DETECT(
        \DB_DETECT[0][29] ), .SB_CORRECT(\SB_CORRECT[0][29] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][29] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[29]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[29]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%7%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C7 (.A_DOUT({
        nc897, nc898, nc899, nc900, nc901, nc902, nc903, nc904, nc905, 
        nc906, nc907, nc908, nc909, nc910, nc911, nc912, nc913, nc914, 
        nc915, R_DATA[7]}), .B_DOUT({nc916, nc917, nc918, nc919, nc920, 
        nc921, nc922, nc923, nc924, nc925, nc926, nc927, nc928, nc929, 
        nc930, nc931, nc932, nc933, nc934, nc935}), .DB_DETECT(
        \DB_DETECT[0][7] ), .SB_CORRECT(\SB_CORRECT[0][7] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][7] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[7]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[7]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%14%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C14 (.A_DOUT({
        nc936, nc937, nc938, nc939, nc940, nc941, nc942, nc943, nc944, 
        nc945, nc946, nc947, nc948, nc949, nc950, nc951, nc952, nc953, 
        nc954, R_DATA[14]}), .B_DOUT({nc955, nc956, nc957, nc958, 
        nc959, nc960, nc961, nc962, nc963, nc964, nc965, nc966, nc967, 
        nc968, nc969, nc970, nc971, nc972, nc973, nc974}), .DB_DETECT(
        \DB_DETECT[0][14] ), .SB_CORRECT(\SB_CORRECT[0][14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][14] ), .A_ADDR({R_ADDR[13], 
        R_ADDR[12], R_ADDR[11], R_ADDR[10], R_ADDR[9], R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0]}), .A_BLK_EN({VCC, VCC, VCC}), 
        .A_CLK(CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND}), 
        .A_REN(R_EN), .A_WEN({GND, GND}), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({W_ADDR[13], 
        W_ADDR[12], W_ADDR[11], W_ADDR[10], W_ADDR[9], W_ADDR[8], 
        W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], W_ADDR[3], 
        W_ADDR[2], W_ADDR[1], W_ADDR[0]}), .B_BLK_EN({W_EN, VCC, VCC}), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        W_DATA[14]}), .B_REN(VCC), .B_WEN({GND, WBYTE_EN[14]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, GND, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, GND, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%12%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C12 (.A_DOUT({
        nc975, nc976, nc977, nc978, nc979, nc980, nc981, nc982, nc983, 
        nc984, nc985, nc986, nc987, nc988, nc989, nc990, nc991, nc992, 
        nc993, R_DATA[12]}), .B_DOUT({nc994, nc995, nc996, nc997, 
        nc998, nc999, nc1000, nc1001, nc1002, nc1003, nc1004, nc1005, 
        nc1006, nc1007, nc1008, nc1009, nc1010, nc1011, nc1012, nc1013})
        , .DB_DETECT(\DB_DETECT[0][12] ), .SB_CORRECT(
        \SB_CORRECT[0][12] ), .ACCESS_BUSY(\ACCESS_BUSY[0][12] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[12]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[12]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%13%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C13 (.A_DOUT({
        nc1014, nc1015, nc1016, nc1017, nc1018, nc1019, nc1020, nc1021, 
        nc1022, nc1023, nc1024, nc1025, nc1026, nc1027, nc1028, nc1029, 
        nc1030, nc1031, nc1032, R_DATA[13]}), .B_DOUT({nc1033, nc1034, 
        nc1035, nc1036, nc1037, nc1038, nc1039, nc1040, nc1041, nc1042, 
        nc1043, nc1044, nc1045, nc1046, nc1047, nc1048, nc1049, nc1050, 
        nc1051, nc1052}), .DB_DETECT(\DB_DETECT[0][13] ), .SB_CORRECT(
        \SB_CORRECT[0][13] ), .ACCESS_BUSY(\ACCESS_BUSY[0][13] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[13]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[13]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%11%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C11 (.A_DOUT({
        nc1053, nc1054, nc1055, nc1056, nc1057, nc1058, nc1059, nc1060, 
        nc1061, nc1062, nc1063, nc1064, nc1065, nc1066, nc1067, nc1068, 
        nc1069, nc1070, nc1071, R_DATA[11]}), .B_DOUT({nc1072, nc1073, 
        nc1074, nc1075, nc1076, nc1077, nc1078, nc1079, nc1080, nc1081, 
        nc1082, nc1083, nc1084, nc1085, nc1086, nc1087, nc1088, nc1089, 
        nc1090, nc1091}), .DB_DETECT(\DB_DETECT[0][11] ), .SB_CORRECT(
        \SB_CORRECT[0][11] ), .ACCESS_BUSY(\ACCESS_BUSY[0][11] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[11]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[11]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%3%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C3 (.A_DOUT({
        nc1092, nc1093, nc1094, nc1095, nc1096, nc1097, nc1098, nc1099, 
        nc1100, nc1101, nc1102, nc1103, nc1104, nc1105, nc1106, nc1107, 
        nc1108, nc1109, nc1110, R_DATA[3]}), .B_DOUT({nc1111, nc1112, 
        nc1113, nc1114, nc1115, nc1116, nc1117, nc1118, nc1119, nc1120, 
        nc1121, nc1122, nc1123, nc1124, nc1125, nc1126, nc1127, nc1128, 
        nc1129, nc1130}), .DB_DETECT(\DB_DETECT[0][3] ), .SB_CORRECT(
        \SB_CORRECT[0][3] ), .ACCESS_BUSY(\ACCESS_BUSY[0][3] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[3]}), .B_REN(VCC), .B_WEN({GND, 
        WBYTE_EN[3]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%30%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C30 (.A_DOUT({
        nc1131, nc1132, nc1133, nc1134, nc1135, nc1136, nc1137, nc1138, 
        nc1139, nc1140, nc1141, nc1142, nc1143, nc1144, nc1145, nc1146, 
        nc1147, nc1148, nc1149, R_DATA[30]}), .B_DOUT({nc1150, nc1151, 
        nc1152, nc1153, nc1154, nc1155, nc1156, nc1157, nc1158, nc1159, 
        nc1160, nc1161, nc1162, nc1163, nc1164, nc1165, nc1166, nc1167, 
        nc1168, nc1169}), .DB_DETECT(\DB_DETECT[0][30] ), .SB_CORRECT(
        \SB_CORRECT[0][30] ), .ACCESS_BUSY(\ACCESS_BUSY[0][30] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[30]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[30]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%2%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C2 (.A_DOUT({
        nc1170, nc1171, nc1172, nc1173, nc1174, nc1175, nc1176, nc1177, 
        nc1178, nc1179, nc1180, nc1181, nc1182, nc1183, nc1184, nc1185, 
        nc1186, nc1187, nc1188, R_DATA[2]}), .B_DOUT({nc1189, nc1190, 
        nc1191, nc1192, nc1193, nc1194, nc1195, nc1196, nc1197, nc1198, 
        nc1199, nc1200, nc1201, nc1202, nc1203, nc1204, nc1205, nc1206, 
        nc1207, nc1208}), .DB_DETECT(\DB_DETECT[0][2] ), .SB_CORRECT(
        \SB_CORRECT[0][2] ), .ACCESS_BUSY(\ACCESS_BUSY[0][2] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[2]}), .B_REN(VCC), .B_WEN({GND, 
        WBYTE_EN[2]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%20%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C20 (.A_DOUT({
        nc1209, nc1210, nc1211, nc1212, nc1213, nc1214, nc1215, nc1216, 
        nc1217, nc1218, nc1219, nc1220, nc1221, nc1222, nc1223, nc1224, 
        nc1225, nc1226, nc1227, R_DATA[20]}), .B_DOUT({nc1228, nc1229, 
        nc1230, nc1231, nc1232, nc1233, nc1234, nc1235, nc1236, nc1237, 
        nc1238, nc1239, nc1240, nc1241, nc1242, nc1243, nc1244, nc1245, 
        nc1246, nc1247}), .DB_DETECT(\DB_DETECT[0][20] ), .SB_CORRECT(
        \SB_CORRECT[0][20] ), .ACCESS_BUSY(\ACCESS_BUSY[0][20] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[20]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[20]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%6%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C6 (.A_DOUT({
        nc1248, nc1249, nc1250, nc1251, nc1252, nc1253, nc1254, nc1255, 
        nc1256, nc1257, nc1258, nc1259, nc1260, nc1261, nc1262, nc1263, 
        nc1264, nc1265, nc1266, R_DATA[6]}), .B_DOUT({nc1267, nc1268, 
        nc1269, nc1270, nc1271, nc1272, nc1273, nc1274, nc1275, nc1276, 
        nc1277, nc1278, nc1279, nc1280, nc1281, nc1282, nc1283, nc1284, 
        nc1285, nc1286}), .DB_DETECT(\DB_DETECT[0][6] ), .SB_CORRECT(
        \SB_CORRECT[0][6] ), .ACCESS_BUSY(\ACCESS_BUSY[0][6] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[6]}), .B_REN(VCC), .B_WEN({GND, 
        WBYTE_EN[6]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%38%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C38 (.A_DOUT({
        nc1287, nc1288, nc1289, nc1290, nc1291, nc1292, nc1293, nc1294, 
        nc1295, nc1296, nc1297, nc1298, nc1299, nc1300, nc1301, nc1302, 
        nc1303, nc1304, nc1305, R_DATA[38]}), .B_DOUT({nc1306, nc1307, 
        nc1308, nc1309, nc1310, nc1311, nc1312, nc1313, nc1314, nc1315, 
        nc1316, nc1317, nc1318, nc1319, nc1320, nc1321, nc1322, nc1323, 
        nc1324, nc1325}), .DB_DETECT(\DB_DETECT[0][38] ), .SB_CORRECT(
        \SB_CORRECT[0][38] ), .ACCESS_BUSY(\ACCESS_BUSY[0][38] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[38]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[38]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%36%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C36 (.A_DOUT({
        nc1326, nc1327, nc1328, nc1329, nc1330, nc1331, nc1332, nc1333, 
        nc1334, nc1335, nc1336, nc1337, nc1338, nc1339, nc1340, nc1341, 
        nc1342, nc1343, nc1344, R_DATA[36]}), .B_DOUT({nc1345, nc1346, 
        nc1347, nc1348, nc1349, nc1350, nc1351, nc1352, nc1353, nc1354, 
        nc1355, nc1356, nc1357, nc1358, nc1359, nc1360, nc1361, nc1362, 
        nc1363, nc1364}), .DB_DETECT(\DB_DETECT[0][36] ), .SB_CORRECT(
        \SB_CORRECT[0][36] ), .ACCESS_BUSY(\ACCESS_BUSY[0][36] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[36]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[36]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%28%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C28 (.A_DOUT({
        nc1365, nc1366, nc1367, nc1368, nc1369, nc1370, nc1371, nc1372, 
        nc1373, nc1374, nc1375, nc1376, nc1377, nc1378, nc1379, nc1380, 
        nc1381, nc1382, nc1383, R_DATA[28]}), .B_DOUT({nc1384, nc1385, 
        nc1386, nc1387, nc1388, nc1389, nc1390, nc1391, nc1392, nc1393, 
        nc1394, nc1395, nc1396, nc1397, nc1398, nc1399, nc1400, nc1401, 
        nc1402, nc1403}), .DB_DETECT(\DB_DETECT[0][28] ), .SB_CORRECT(
        \SB_CORRECT[0][28] ), .ACCESS_BUSY(\ACCESS_BUSY[0][28] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[28]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[28]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%26%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C26 (.A_DOUT({
        nc1404, nc1405, nc1406, nc1407, nc1408, nc1409, nc1410, nc1411, 
        nc1412, nc1413, nc1414, nc1415, nc1416, nc1417, nc1418, nc1419, 
        nc1420, nc1421, nc1422, R_DATA[26]}), .B_DOUT({nc1423, nc1424, 
        nc1425, nc1426, nc1427, nc1428, nc1429, nc1430, nc1431, nc1432, 
        nc1433, nc1434, nc1435, nc1436, nc1437, nc1438, nc1439, nc1440, 
        nc1441, nc1442}), .DB_DETECT(\DB_DETECT[0][26] ), .SB_CORRECT(
        \SB_CORRECT[0][26] ), .ACCESS_BUSY(\ACCESS_BUSY[0][26] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[26]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[26]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%35%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C35 (.A_DOUT({
        nc1443, nc1444, nc1445, nc1446, nc1447, nc1448, nc1449, nc1450, 
        nc1451, nc1452, nc1453, nc1454, nc1455, nc1456, nc1457, nc1458, 
        nc1459, nc1460, nc1461, R_DATA[35]}), .B_DOUT({nc1462, nc1463, 
        nc1464, nc1465, nc1466, nc1467, nc1468, nc1469, nc1470, nc1471, 
        nc1472, nc1473, nc1474, nc1475, nc1476, nc1477, nc1478, nc1479, 
        nc1480, nc1481}), .DB_DETECT(\DB_DETECT[0][35] ), .SB_CORRECT(
        \SB_CORRECT[0][35] ), .ACCESS_BUSY(\ACCESS_BUSY[0][35] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[35]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[35]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%25%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C25 (.A_DOUT({
        nc1482, nc1483, nc1484, nc1485, nc1486, nc1487, nc1488, nc1489, 
        nc1490, nc1491, nc1492, nc1493, nc1494, nc1495, nc1496, nc1497, 
        nc1498, nc1499, nc1500, R_DATA[25]}), .B_DOUT({nc1501, nc1502, 
        nc1503, nc1504, nc1505, nc1506, nc1507, nc1508, nc1509, nc1510, 
        nc1511, nc1512, nc1513, nc1514, nc1515, nc1516, nc1517, nc1518, 
        nc1519, nc1520}), .DB_DETECT(\DB_DETECT[0][25] ), .SB_CORRECT(
        \SB_CORRECT[0][25] ), .ACCESS_BUSY(\ACCESS_BUSY[0][25] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[25]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[25]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("LSRAM_code%16384-16384%40-40%SPEED%0%17%TWO-PORT")
         )  LSRAM_code_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C17 (.A_DOUT({
        nc1521, nc1522, nc1523, nc1524, nc1525, nc1526, nc1527, nc1528, 
        nc1529, nc1530, nc1531, nc1532, nc1533, nc1534, nc1535, nc1536, 
        nc1537, nc1538, nc1539, R_DATA[17]}), .B_DOUT({nc1540, nc1541, 
        nc1542, nc1543, nc1544, nc1545, nc1546, nc1547, nc1548, nc1549, 
        nc1550, nc1551, nc1552, nc1553, nc1554, nc1555, nc1556, nc1557, 
        nc1558, nc1559}), .DB_DETECT(\DB_DETECT[0][17] ), .SB_CORRECT(
        \SB_CORRECT[0][17] ), .ACCESS_BUSY(\ACCESS_BUSY[0][17] ), 
        .A_ADDR({R_ADDR[13], R_ADDR[12], R_ADDR[11], R_ADDR[10], 
        R_ADDR[9], R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], 
        R_ADDR[4], R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0]}), 
        .A_BLK_EN({VCC, VCC, VCC}), .A_CLK(CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .A_REN(R_EN), .A_WEN({GND, GND}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[13], W_ADDR[12], W_ADDR[11], W_ADDR[10], 
        W_ADDR[9], W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0]}), 
        .B_BLK_EN({W_EN, VCC, VCC}), .B_CLK(CLK), .B_DIN({GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, W_DATA[17]}), .B_REN(VCC), .B_WEN({
        GND, WBYTE_EN[17]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(GND), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, GND, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, GND, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
