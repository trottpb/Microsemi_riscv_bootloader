//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Fri Aug 03 11:38:46 2018
// Version: PolarFire v2.2 12.200.30.10
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// RCOSC
module RCOSC(
    // Outputs
    RCOSC_160MHZ_GL
);

//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output RCOSC_160MHZ_GL;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   RCOSC_160MHZ_GL_0;
wire   RCOSC_160MHZ_GL_0_net_0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign RCOSC_160MHZ_GL_0_net_0 = RCOSC_160MHZ_GL_0;
assign RCOSC_160MHZ_GL         = RCOSC_160MHZ_GL_0_net_0;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------RCOSC_RCOSC_0_PF_OSC   -   Actel:SgCore:PF_OSC:1.0.102
RCOSC_RCOSC_0_PF_OSC RCOSC_0(
        // Outputs
        .RCOSC_160MHZ_GL ( RCOSC_160MHZ_GL_0 ) 
        );


endmodule
